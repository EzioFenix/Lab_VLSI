LIBRARY IEEE;
USE IEEE.Std_logic_1164.ALL;
ENTITY Gen25MHz IS
	PORT (
		clk50MHz : IN STD_LOGIC;
		clk25MHz : INOUT STD_LOGIC := '0');
END ENTITY;
ARCHITECTURE behavior OF Gen25MHZ IS
BEGIN
	PROCESS (clk50MHz)
	BEGIN
		IF clk50MHz'event AND clk50MHz = '1' THEN
			clk25MHz <= NOT clk25MHz;
		END IF;
	END PROCESS;
END behavior;